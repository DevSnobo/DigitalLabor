`timescale 1 ns / 100 ps
module  test_LPM_MULT_20_20_40_SIGNED_1_UNUSED (Result, DataA, DataB,
        Clock, Aclr); // synthesis syn_black_box

input   Clock, Aclr;
input   [19:0]  DataA;
input   [19:0]  DataB;
output  [39:0]  Result;


endmodule

