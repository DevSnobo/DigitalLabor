`timescale 1 ns / 100 ps
module  test (Result, DataA_, DataB_); // synthesis syn_black_box

input   [15:0]  DataA_;
input   [15:0]  DataB_;
output  [31:0]  Result;


endmodule

