module logic12(d1,a2,a3);

input a2,a3;
output d1;

assign d1 = a2 & a3;

endmodule

