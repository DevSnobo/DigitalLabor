module user_nor2(d0,a0,a1);

input a0,a1;
output d0;

assign d0 = !(a0|a1);

endmodule

