library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity test_ent is

end;

architecture test_arch of test_ent is
begin

end test_arch;

